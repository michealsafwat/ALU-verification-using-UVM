package test_pkg;
`include "ALU_IF.svh"
import uvm_pkg::*;
`include "uvm_macros.svh"

  `include "transaction.svh"
  `include "base_sequence.svh"
  `include "sequencer.svh"
  `include "driver.svh"
  `include "monitor.svh"
  `include "coverage.svh"
  `include "scoreboard.svh"
  `include "agent.svh"
  `include "environment.svh"
  `include "test.svh"
endpackage : test_pkg
